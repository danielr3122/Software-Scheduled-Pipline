-------------------------------------------------------------------------
-- Brayton Rude
-- rude87@iastate.edu
-------------------------------------------------------------------------
-- decoder5t32.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 5:32bit decoder.
--
-- 09/22/2022 by BR::Design created.
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity decoder5t32 is
    port(i_A   : in std_logic_vector(4 downto 0);
         o_F   : out std_logic_vector(31 downto 0));
end decoder5t32;

architecture dataflow of decoder5t32 is

begin

    with i_A select
        o_F <=  x"0000_0001" when "00000", -- $0
                x"0000_0002" when "00001", -- $1
                x"0000_0004" when "00010", -- $2
                x"0000_0008" when "00011", -- $3
                x"0000_0010" when "00100", -- $4
                x"0000_0020" when "00101", -- $5
                x"0000_0040" when "00110", -- $6
                x"0000_0080" when "00111", -- $7
                x"0000_0100" when "01000", -- $8
                x"0000_0200" when "01001", -- $9
                x"0000_0400" when "01010", -- $10
                x"0000_0800" when "01011", -- $11
                x"0000_1000" when "01100", -- $12
                x"0000_2000" when "01101", -- $13
                x"0000_4000" when "01110", -- $14
                x"0000_8000" when "01111", -- $15
                x"0001_0000" when "10000", -- $16
                x"0002_0000" when "10001", -- $17
                x"0004_0000" when "10010", -- $18
                x"0008_0000" when "10011", -- $19
                x"0010_0000" when "10100", -- $20
                x"0020_0000" when "10101", -- $21
                x"0040_0000" when "10110", -- $22
                x"0080_0000" when "10111", -- $23
                x"0100_0000" when "11000", -- $24
                x"0200_0000" when "11001", -- $25
                x"0400_0000" when "11010", -- $26
                x"0800_0000" when "11011", -- $27
                x"1000_0000" when "11100", -- $28
                x"2000_0000" when "11101", -- $29
                x"4000_0000" when "11110", -- $30
                x"8000_0000" when "11111", -- $31
                x"0000_0000" when others;  -- Error

end dataflow;